library verilog;
use verilog.vl_types.all;
entity tb_core_ut is
end tb_core_ut;
