library verilog;
use verilog.vl_types.all;
entity rv32_assembler is
end rv32_assembler;
