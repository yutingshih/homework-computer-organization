library verilog;
use verilog.vl_types.all;
entity kronos_types is
end kronos_types;
