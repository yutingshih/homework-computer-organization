library verilog;
use verilog.vl_types.all;
entity reg00 is
    port(
        x0              : in     vl_logic_vector(31 downto 0);
        x1              : in     vl_logic_vector(31 downto 0);
        x2              : in     vl_logic_vector(31 downto 0);
        x3              : in     vl_logic_vector(31 downto 0);
        x4              : in     vl_logic_vector(31 downto 0);
        x5              : in     vl_logic_vector(31 downto 0);
        x6              : in     vl_logic_vector(31 downto 0);
        x7              : in     vl_logic_vector(31 downto 0);
        x8              : in     vl_logic_vector(31 downto 0);
        x9              : in     vl_logic_vector(31 downto 0);
        x10             : in     vl_logic_vector(31 downto 0);
        x11             : in     vl_logic_vector(31 downto 0);
        x12             : in     vl_logic_vector(31 downto 0);
        x13             : in     vl_logic_vector(31 downto 0);
        x14             : in     vl_logic_vector(31 downto 0);
        x15             : in     vl_logic_vector(31 downto 0);
        x16             : in     vl_logic_vector(31 downto 0);
        x17             : in     vl_logic_vector(31 downto 0);
        x18             : in     vl_logic_vector(31 downto 0);
        x19             : in     vl_logic_vector(31 downto 0);
        x20             : in     vl_logic_vector(31 downto 0);
        x21             : in     vl_logic_vector(31 downto 0);
        x22             : in     vl_logic_vector(31 downto 0);
        x23             : in     vl_logic_vector(31 downto 0);
        x24             : in     vl_logic_vector(31 downto 0);
        x25             : in     vl_logic_vector(31 downto 0);
        x26             : in     vl_logic_vector(31 downto 0);
        x27             : in     vl_logic_vector(31 downto 0);
        x28             : in     vl_logic_vector(31 downto 0);
        x29             : in     vl_logic_vector(31 downto 0);
        x30             : in     vl_logic_vector(31 downto 0);
        x31             : in     vl_logic_vector(31 downto 0)
    );
end reg00;
